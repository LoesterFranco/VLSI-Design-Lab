*LAB - 5 - Studythe behaviour transfer function, Noise margin, effect on risetime, falltime, propagation delay, power and energy consumec of CMOS gates like NAND, NOR, functions like AOI and 2 input XOR gate with variation in L and W of the pullup and pulldown transistors. Also power consumed with non ideal step input. Study the effect of VSB due to series connected transistors.

.include ./level3.txt

* 3 input AOI GATE

mpa nabc a pos pos cmosp w=4u l=1u
mpb nabc b pos pos cmosp w=4u l=1u
mpb out c nabc pos cmosp w=4u l=1u
mna out a nab 0 cmosn w=1u l=1u
mnb nab b 0 0 cmosn w=1u l=1u 
mnc out c 0 0 cmosn w=1u l=1u 

*vout1 out out1 0
*vout2 out out2 0
vpos pos 0 5
va a 0 0 pulse(0 5 4n 0.1n 0.1n 3.8n 8n)
vb b 0 0 pulse(0 5 2n 0.1n 0.1n 1.8n 4n)

vc c 0 0 pulse(0 5 1n 0.1n 0.1n 0.8n 2n)


.control
		tran 0.01n 8n
		plot v(a) v(b) v(c) v(out)
		let power = -5*vpos#branch
		meas tran pavg AVG power from=0n to=4n
.endc
.end

