magic
tech scmos
timestamp 1603383315
<< polysilicon >>
rect 31 51 33 53
rect 31 37 33 42
rect -12 35 33 37
rect -12 6 -10 35
rect 31 32 33 35
rect 31 27 33 29
rect 25 21 87 23
rect 25 6 27 21
rect -9 3 -8 5
rect 1 3 3 5
rect 12 3 14 5
rect 23 3 24 5
rect -12 -19 -10 2
rect 85 5 87 21
rect 51 3 52 5
rect 61 3 63 5
rect 72 3 74 5
rect 83 3 87 5
rect -12 -21 -5 -19
rect -2 -21 0 -19
rect 25 -20 27 2
rect 8 -22 10 -20
rect 13 -22 27 -20
rect 48 -19 50 2
rect 48 -21 55 -19
rect 58 -21 60 -19
rect 85 -20 87 3
rect 96 19 170 21
rect 96 -7 98 19
rect 108 3 112 5
rect 121 3 123 5
rect 132 3 134 5
rect 143 3 144 5
rect 68 -22 70 -20
rect 73 -22 87 -20
rect 108 -19 110 3
rect 168 5 170 19
rect 168 3 172 5
rect 181 3 183 5
rect 192 3 194 5
rect 203 3 207 5
rect 108 -21 115 -19
rect 118 -21 120 -19
rect 145 -20 147 2
rect 108 -40 110 -21
rect 128 -22 130 -20
rect 133 -22 147 -20
rect 154 -32 156 -11
rect 168 -19 170 3
rect 168 -21 175 -19
rect 178 -21 180 -19
rect 205 -20 207 3
rect 188 -22 190 -20
rect 193 -22 207 -20
rect 205 -32 207 -22
rect 154 -34 207 -32
rect 102 -42 110 -40
<< ndiffusion >>
rect 29 29 31 32
rect 33 29 35 32
rect -5 -19 -2 -17
rect 10 -20 13 -18
rect -5 -23 -2 -21
rect 55 -19 58 -17
rect 70 -20 73 -18
rect 10 -24 13 -22
rect 55 -23 58 -21
rect 115 -19 118 -17
rect 130 -20 133 -18
rect 70 -24 73 -22
rect 115 -23 118 -21
rect 130 -24 133 -22
rect 175 -19 178 -17
rect 190 -20 193 -18
rect 175 -23 178 -21
rect 190 -24 193 -22
<< pdiffusion >>
rect 28 49 31 51
rect 29 45 31 49
rect 28 42 31 45
rect 33 49 36 51
rect 33 45 35 49
rect 33 42 36 45
rect -8 7 -6 8
rect -2 7 1 8
rect -8 5 1 7
rect 14 7 16 8
rect 20 7 23 8
rect 14 5 23 7
rect 52 7 54 8
rect 58 7 61 8
rect -8 1 1 3
rect -8 0 -6 1
rect -2 0 1 1
rect 14 1 23 3
rect 52 5 61 7
rect 74 7 76 8
rect 80 7 83 8
rect 74 5 83 7
rect 14 0 16 1
rect 20 0 23 1
rect 52 1 61 3
rect 52 0 54 1
rect 58 0 61 1
rect 74 1 83 3
rect 74 0 76 1
rect 80 0 83 1
rect 112 7 114 8
rect 118 7 121 8
rect 112 5 121 7
rect 134 7 136 8
rect 140 7 143 8
rect 134 5 143 7
rect 112 1 121 3
rect 112 0 114 1
rect 118 0 121 1
rect 134 1 143 3
rect 172 7 174 8
rect 178 7 181 8
rect 172 5 181 7
rect 194 7 196 8
rect 200 7 203 8
rect 194 5 203 7
rect 134 0 136 1
rect 140 0 143 1
rect 172 1 181 3
rect 172 0 174 1
rect 178 0 181 1
rect 194 1 203 3
rect 194 0 196 1
rect 200 0 203 1
<< metal1 >>
rect 20 54 66 58
rect 20 49 24 54
rect 10 45 25 49
rect 10 15 14 45
rect 39 39 43 49
rect 39 35 51 39
rect 39 28 43 35
rect 25 21 29 28
rect 25 17 36 21
rect -6 11 20 15
rect -6 -7 -2 -3
rect 16 -7 20 -3
rect -21 -11 20 -7
rect -21 -39 -17 -11
rect -6 -13 -2 -11
rect 2 -18 9 -14
rect 2 -23 6 -18
rect -2 -27 6 -23
rect 32 -24 36 17
rect 47 6 51 35
rect 62 15 66 54
rect 54 11 200 15
rect 148 2 166 6
rect 54 -7 58 -3
rect 76 -7 80 -3
rect 114 -7 118 -3
rect 136 -7 140 -3
rect 162 -7 166 2
rect 174 -7 178 -3
rect 196 -7 200 -3
rect 54 -11 95 -7
rect 114 -11 153 -7
rect 162 -11 200 -7
rect 54 -13 58 -11
rect 114 -13 118 -11
rect 62 -18 69 -14
rect 174 -13 178 -11
rect 122 -18 129 -14
rect 182 -18 189 -14
rect 62 -23 66 -18
rect 122 -23 126 -18
rect 182 -23 186 -18
rect 13 -28 36 -24
rect 58 -27 66 -23
rect 32 -31 36 -28
rect 118 -27 126 -23
rect 69 -31 73 -28
rect 178 -27 186 -23
rect 129 -31 133 -28
rect 189 -31 193 -28
rect 32 -35 193 -31
rect -21 -43 98 -39
<< ntransistor >>
rect 31 29 33 32
rect -5 -21 -2 -19
rect 10 -22 13 -20
rect 55 -21 58 -19
rect 70 -22 73 -20
rect 115 -21 118 -19
rect 130 -22 133 -20
rect 175 -21 178 -19
rect 190 -22 193 -20
<< ptransistor >>
rect 31 42 33 51
rect -8 3 1 5
rect 14 3 23 5
rect 52 3 61 5
rect 74 3 83 5
rect 112 3 121 5
rect 134 3 143 5
rect 172 3 181 5
rect 194 3 203 5
<< polycontact >>
rect -13 2 -9 6
rect 24 2 28 6
rect 47 2 51 6
rect 95 -11 99 -7
rect 144 2 148 6
rect 153 -11 157 -7
rect 98 -43 102 -39
<< ndcontact >>
rect 25 28 29 32
rect 35 28 39 32
rect -6 -17 -2 -13
rect 9 -18 13 -14
rect 54 -17 58 -13
rect 69 -18 73 -14
rect -6 -27 -2 -23
rect 114 -17 118 -13
rect 129 -18 133 -14
rect 9 -28 13 -24
rect 54 -27 58 -23
rect 69 -28 73 -24
rect 114 -27 118 -23
rect 129 -28 133 -24
rect 174 -17 178 -13
rect 189 -18 193 -14
rect 174 -27 178 -23
rect 189 -28 193 -24
<< pdcontact >>
rect 25 45 29 49
rect 35 45 39 49
rect -6 7 -2 11
rect 16 7 20 11
rect 54 7 58 11
rect -6 -3 -2 1
rect 76 7 80 11
rect 16 -3 20 1
rect 54 -3 58 1
rect 76 -3 80 1
rect 114 7 118 11
rect 136 7 140 11
rect 114 -3 118 1
rect 174 7 178 11
rect 196 7 200 11
rect 136 -3 140 1
rect 174 -3 178 1
rect 196 -3 200 1
<< labels >>
rlabel polycontact -11 4 -11 4 1 D
rlabel metal1 42 56 42 56 5 Vdd
rlabel polycontact 26 4 26 4 1 clock
rlabel metal1 92 -33 92 -33 1 0
rlabel polycontact 49 4 49 4 1 Dbar
rlabel polycontact 100 -41 100 -41 1 S
rlabel polycontact 97 -9 97 -9 1 R
rlabel polycontact 155 -9 155 -9 1 Q
rlabel polycontact 146 4 146 4 1 Qbar
<< end >>
