magic
tech scmos
timestamp 242945690
<< polysilicon >>
rect -13 15 -11 17
rect 3 15 5 17
rect -13 6 -11 9
rect -14 2 -11 6
rect 3 5 5 9
rect -13 -1 -11 2
rect -2 3 5 5
rect 3 -1 5 3
rect -13 -9 -11 -7
rect 3 -9 5 -7
<< ndiffusion >>
rect -16 -2 -13 -1
rect -14 -6 -13 -2
rect -16 -7 -13 -6
rect -11 -2 -8 -1
rect 0 -2 3 -1
rect -11 -6 -10 -2
rect 2 -6 3 -2
rect -11 -7 -8 -6
rect 0 -7 3 -6
rect 5 -2 8 -1
rect 5 -6 6 -2
rect 5 -7 9 -6
<< pdiffusion >>
rect -16 14 -13 15
rect -14 10 -13 14
rect -16 9 -13 10
rect -11 14 -8 15
rect 0 14 3 15
rect -11 10 -10 14
rect 2 10 3 14
rect -11 9 -8 10
rect 0 9 3 10
rect 5 14 8 15
rect 5 10 6 14
rect 5 9 8 10
<< metal1 >>
rect -9 18 10 21
rect -18 14 -15 17
rect -9 14 -6 18
rect 7 14 10 18
rect -3 10 -2 13
rect -3 8 0 10
rect 7 -2 10 10
91rect -6 -6 -2 -3
rect -18 -8 -15 -6
<< ntransistor >>
rect -13 -7 -11 -1
rect 3 -7 5 -1
<< ptransistor >>
rect -13 9 -11 15
rect 3 9 5 15
<< polycontact >>
rect -18 2 -14 6
rect -6 1 -2 5
<< ndcontact >>
rect -18 -6 -14 -2
rect -10 -6 -6 -2
rect -2 -6 2 -2
rect 6 -6 10 -2
<< pdcontact >>
rect -18 10 -14 14
rect -10 10 -6 14
rect -2 10 2 14
rect 6 10 10 14
<< labels >>
rlabel metal1 -17 16 -17 16 5 vdd
rlabel metal1 9 4 9 4 5 out
rlabel polycontact -4 3 -4 3 5 in2
rlabel polycontact -16 4 -16 4 5 in1
rlabel metal1 -17 -7 -17 -7 3 0
rlabel metal1 -4 -5 -4 -5 1 x
rlabel metal1 -2 9 -2 9 5 vdd
<< end >>