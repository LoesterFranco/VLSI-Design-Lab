magic
tech scmos
timestamp 2602923583
<< polysilicon >>
rect -1 18 1 20
rect 10 19 25 21
rect 15 18 17 19
rect -1 3 1 6
rect 15 4 17 6
rect -2 -1 1 3
rect -1 -4 1 -1
rect 15 -4 17 -2
rect -1 -9 1 -7
rect 15 -10 17 -7
rect 23 -10 25 19
rect 15 -12 25 -10
<< ndiffusion >>
rect -2 -7 -1 -4
rect 1 -7 2 -4
rect 14 -7 15 -4
rect 17 -7 18 -4
<< pdiffusion >>
rect -4 11 -1 18
rect -2 7 -1 11
rect -4 6 -1 7
rect 1 11 4 18
rect 12 11 15 18
rect 1 7 2 11
rect 14 7 15 11
rect 1 6 4 7
rect 12 6 15 7
rect 17 11 20 18
rect 17 7 18 11
rect 17 6 20 7
<< metal1 >>
rect -6 11 -3 20
rect 6 7 10 10
rect 19 2 22 7
rect 3 -1 22 2
rect 3 -4 6 -1
rect 19 -4 22 -1
rect -6 -11 -3 -8
rect 11 -11 14 -8
rect -6 -14 14 -11
<< ntransistor >>
rect -1 -7 1 -4
rect 15 -7 17 -4
<< ptransistor >>
rect -1 6 1 18
rect 15 6 17 18
<< polycontact >>
rect 6 17 10 21
rect -6 -1 -2 3
<< ndcontact >>
rect -6 -8 -2 -4
rect 2 -8 6 -4
rect 10 -8 14 -4
rect 18 -8 22 -4
<< pdcontact >>
rect -6 7 -2 11
rect 2 7 6 11
rect 10 7 14 11
rect 18 7 22 11
<< labels >>
rlabel metal1 -5 19 -5 19 5 vdd
rlabel metal1 8 1 8 1 5 out
rlabel metal1 8 9 8 9 5 x
rlabel polycontact 8 19 8 19 1 in2
rlabel polycontact -4 1 -4 1 1 in1
rlabel metal1 4 -13 4 -13 1 0
<< end >>